module MIPS_Cpu_Control #(
    parameters
    //take in op code (31-26)
)
//figure out what command the opcode corresponds to

//set RegDst, ALUSRC, MemtoReg, RegWrite, MemRead, MemWrite, Branch, ALUOp1, ALUOp0
//to their correspoding bits

//Use switch statement most likely

//ex
//if instruction is lw
    //RegDst = 0
    //ALUSrc = 1
    //MemtoReg = 1
    //etc...

//if jump, composition is different


endmodule