module MIPS_Cpu_Core #(
    parameters
)


endmodule