module MIPS_Cpu_Top #(
    parameters
)

MIPS_Cpu_Control cpu_cont (

)

endmodule