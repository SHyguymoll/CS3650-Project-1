module MIPS_Cpu_Top #(
    parameters
)
    //Pass the instruction into control to get the signals
    //Pass the signal effects along with rest of instructions into core
    
MIPS_Cpu_Control cpu_cont (

)

endmodule