module MIPS_Cpu_Control #(
    parameters
)



endmodule